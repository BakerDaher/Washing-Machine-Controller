LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SevSeg_Decoder IS
 PORT ( INPUT : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		  SEVSEG_BUS : OUT STD_LOGIC_VECTOR (6 DOWNTO 0));
END SevSeg_Decoder;

ARCHITECTURE BEHAVIORAL OF SevSeg_Decoder IS

BEGIN

WITH INPUT SELECT SEVSEG_BUS <=
"1111110" WHEN "00000", --0
"0110000" WHEN "00001", --1
"1101101" WHEN "00010", --2 
"1111001" WHEN "00011", --3 
"0110011" WHEN "00100", --4 
"1011011" WHEN "00101", --5 
"1011111" WHEN "00110", --6 
"1110000" WHEN "00111", --7 
"1111111" WHEN "01000", --8 
"1111011" WHEN "01001", --9 
"1110111" WHEN "01010", --A 
"1111111" WHEN "01011", --B 
"1001110" WHEN "01100", --C 
"1111110" WHEN "01101", --D 
"1001111" WHEN "01110", --E
"0001110" WHEN "01111", --L

"0011110" WHEN "10000", -- W Part left 1
"0111100" WHEN "10001", -- W Part right 2
"1110110" WHEN "10010", -- N 
"1100111" WHEN "10011", -- P
"1100111" WHEN "10100", -- R
"1011011" WHEN "10101", -- S   
"1000011" WHEN "10110", -- T
"0110111" WHEN "10111", -- H
"0000111" WHEN "11000", -- K
"1100111" WHEN "11001", -- P
"0000110" WHEN "11011", -- I 
"1111110" WHEN "11101", -- O
"0000000" WHEN "11010", -- Blank
"0000000" WHEN OTHERS;
END BEHAVIORAL;